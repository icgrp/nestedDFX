module reconfig_inst(
   input rst,
   input gclk,
   output [3:0] upper,
   output [3:0] lower
   );
endmodule
